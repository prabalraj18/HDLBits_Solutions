//Exams/m2014 q4i
module top_module (
    output out);

    assign out = 0 ;
    
endmodule

