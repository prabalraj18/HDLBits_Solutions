// Zero
module top_module(output zero)
    
   assign zero = 1'b0;

endmodule

